module Part1(SW,CLOCK_50,LEDR,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5);
input [9:0] SW;
input CLOCK_50;
output [9:0] LEDR;
output [6:0] HEX0,HEX1,HEX2,HEX3,HEX4,HEX5;





endmodule  